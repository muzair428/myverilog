module full_adders(
    
);
    
endmodule