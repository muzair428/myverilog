module gate2 (
    input wire a,
    input wire b,
    input wire c,
    input wire d,
    input wire e,
    input wire l,

    output wire t,
    output wire k,
);

assign f=(u^j);
assign t=!(e|f);
assign k=!(l&f);
    
endmodule